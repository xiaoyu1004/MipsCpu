`include "cpu.vh"

module ex_stage(
  input                         clk           ,
  input                         reset         ,
  // allouin
  input                         ms_allowin    ,
  output                        es_allowin    ,
  
);
endmodule
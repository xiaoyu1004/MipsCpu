`include "cpu.vh"

module alu(
  input   [11:0]  alu_op    ,
  input   [31:0]  alu_src1  ,
  input   [31:0]  alu_src2  ,
  output  [31:0] alu_result 
);
endmodule